library verilog;
use verilog.vl_types.all;
entity Exp1_vlg_vec_tst is
end Exp1_vlg_vec_tst;
