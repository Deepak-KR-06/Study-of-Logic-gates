library verilog;
use verilog.vl_types.all;
entity Exp1_vlg_check_tst is
    port(
        c               : in     vl_logic;
        d               : in     vl_logic;
        e               : in     vl_logic;
        f               : in     vl_logic;
        g               : in     vl_logic;
        h               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Exp1_vlg_check_tst;
