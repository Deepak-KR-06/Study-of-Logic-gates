library verilog;
use verilog.vl_types.all;
entity Exp1 is
    port(
        a               : in     vl_logic;
        b               : in     vl_logic;
        c               : out    vl_logic;
        d               : out    vl_logic;
        e               : out    vl_logic;
        f               : out    vl_logic;
        g               : out    vl_logic;
        h               : out    vl_logic
    );
end Exp1;
